`default_nettype none

module TuringMachine_test();
  logic [3:0] input_data;
  logic clock, Reset, Next, Done;
  logic [5:0] next_state_out;
  logic [1:0] direction;
  logic [5:0] data_reg_out;

  TuringMachine #(4, 64) dut (.*);

  initial begin
    clock = 1'b0;
    forever #5 clock = ~clock;
  end

  initial begin
    $monitor($time,, "input_data = %d, next = %b, done = %b, next_state_out = %d \
direction = %d, data_reg_out = %d",
             input_data, Next, Done, next_state_out, direction, data_reg_out);
    Reset <= 1'b1;
    Next <= 1'b0; Done <= 1'b0;
    @(posedge clock);
    Reset <= 1'b0;
    input_data <= 3;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 2;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 3;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 2;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 2;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 3;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 3;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 1;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);
    input_data <= 0;
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    @(posedge clock);

    Done <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Done <= 1'b0;
    @(posedge clock);
    @(posedge clock);

    if ((next_state_out != 1) || (direction != 2) || (data_reg_out != 6'b000001)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 1) || (direction != 2) || (data_reg_out != 6'b000011)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 1) || (direction != 2) || (data_reg_out != 6'b000111)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 1) || (direction != 2) || (data_reg_out != 6'b001111)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 2) || (direction != 2) || (data_reg_out != 6'b011110)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 3) || (direction != 1) || (data_reg_out != 6'b111111)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 2) || (direction != 2) || (data_reg_out != 6'b111111)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 2) || (direction != 2) || (data_reg_out != 6'b111111)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 3) || (direction != 1) || (data_reg_out != 6'b111110)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 3) || (direction != 3) || (data_reg_out != 6'b111100)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b1;
    @(posedge clock);
    @(posedge clock);
    Next <= 1'b0;
    @(posedge clock);
    if ((next_state_out != 3) || (direction != 3) || (data_reg_out != 6'b111100)) {
      $$display("next state error\n");
    }
    @(posedge clock);
    #1 $finish;
  end

endmodule: TuringMachine_test